module DW_ecc_width4_chkbits5_synd_sel1(gen, correct_n, datain, chkin,
     err_detect, err_multpl, dataout, chkout);
  input gen, correct_n;
  input [3:0] datain;
  input [4:0] chkin;
  output err_detect, err_multpl;
  output [3:0] dataout;
  output [4:0] chkout;
  wire gen, correct_n;
  wire [3:0] datain;
  wire [4:0] chkin;
  wire err_detect, err_multpl;
  wire [3:0] dataout;
  wire [4:0] chkout;
endmodule