module test #(
    parameter int ROWS = 4,
    parameter int COLS = 8,
    parameter int WIDTH = 16
)(
    input logic [WIDTH-1:0] data_in [ROWS][COLS]
);

endmodule
